version https://git-lfs.github.com/spec/v1
oid sha256:bde83157f82ccb2bb025c704a7837678b708be68c55eb2d09fb973cb08ded229
size 68510854
