version https://git-lfs.github.com/spec/v1
oid sha256:b043de9ce01fac1ef6d7a1bdf7123d5be1db88a415d76d0cd4e2764d94237665
size 170279
